parameter num_of_bits = 1;
